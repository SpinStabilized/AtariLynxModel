* -------------------------------------------------------------------
* 4069 Hex Inverter
* Brian McLaughlin - bjmclaughlin@gmail.com
* -------------------------------------------------------------------
* Connections: A
*              |  Not A
*              |  |  B
*              |  |  |  Not B
*              |  |  |  |
*              |  |  |  |  C
*              |  |  |  |  |  Not C
*              |  |  |  |  |  |  Vss
*              |  |  |  |  |  |  |   Not_D
*              |  |  |  |  |  |  |   |  D
*              |  |  |  |  |  |  |   |  |  Not_E
*              |  |  |  |  |  |  |   |  |  |   E
*              |  |  |  |  |  |  |   |  |  |  |  Not_F
*              |  |  |  |  |  |  |   |  |  |  |  |  F
*              |  |  |  |  |  |  |   |  |  |  |  |  |  Vdd
*              |  |  |  |  |  |  |   |  |  |  |  |  |  |
.SUBCKT 4069IC A  NA B  NB C  NC Vss ND D  NE E  NF F  Vdd

XA A NA Vdd Vss 4069Gate
XB B NB Vdd Vss 4069Gate
XC C NC Vdd Vss 4069Gate
XD D ND Vdd Vss 4069Gate
XE E NE Vdd Vss 4069Gate
XF F NF Vdd Vss 4069Gate

.ENDS 4069IC

* -------------------------------------------------------------------
* 4069 Hex Gate
* -------------------------------------------------------------------
.SUBCKT 4069Gate IN OUT Vdd Vss

M1 IN OUT Vdd Vdd CD4069BP
M2 IN OUT Vss Vss CD4069BN

.MODEL CD4069BN NMOS (LEVEL=1 VTO=2.1 KP=2.9M GAMMA=3.97U
+ PHI=.75 LAMBDA=1.87M RD=20.2 RS=184.1 IS=31.2F PB=.8 MJ=.46
+ CBD=47.6P CBS=57.2P CGSO=70.2N CGDO=58.5N CGBO=96.3N)

.MODEL CD4069BP PMOS (LEVEL=1 VTO=-2.9 KP=2M GAMMA=3.97U
+ PHI=.75 LAMBDA=1.87M RD=28.2 RS=145.2 IS=31.2F PB=.8 MJ=.46
+ CBD=47.6P CBS=57.2P CGSO=70.2N CGDO=58.5N CGBO=96.3N)

.ENDS
* -------------------------------------------------------------------
