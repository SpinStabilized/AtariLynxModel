* -----------------------------------------------------------------------------
* 1N5991B Zener Model - Approximated from Diodes Inc BZT52C4V3
* Brian McLaughlin - bjmclaughlin@gmail.com
*
* Reference: http://www.diodes.com/spicemodels/search.php
*
* Sub-circuit Connections
* A K
* -----------------------------------------------------------------------------
.SUBCKT 1N5991B  A K

.MODEL DF D ( IS=47.9p RS=35.4 N=1.10 CJO=370p VJ=0.750 M=0.330 TT=50.1n )
.MODEL DR D ( IS=9.58f RS=74.5 N=3.00 )

D1 A K DF
DZ 3 A DR
VZ K 3 1.83

.ENDS 1N5991B
