* -----------------------------------------------------------------------------
* SBT-0260 DC Line Filter
* Brian McLaughlin - bjmclaughlin@gmail.com
* -----------------------------------------------------------------------------
.SUBCKT SBT0260 1 2

L1 1 3 60u
R1 3 2 50m

.ENDS SBT0260
